*** SPICE deck for cell 5BitDac_sim_digital{sch} from library Lab_1_DAC
*** Created on Wed Sep 24, 2025 16:22:55
*** Last revised on Wed Sep 24, 2025 16:30:26
*** Written on Wed Sep 24, 2025 16:38:44 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Lab_1_DAC__SingleCell FROM CELL SingleCell{sch}
.SUBCKT Lab_1_DAC__SingleCell bot in out
Rresnwell@0 net@1 in 10k
Rresnwell@1 out net@1 10k
Rresnwell@2 out bot 10k
.ENDS Lab_1_DAC__SingleCell

*** SUBCIRCUIT Lab_1_DAC__5BitDAC FROM CELL 5BitDAC{sch}
.SUBCKT Lab_1_DAC__5BitDAC b0 b1 b2 b3 b4 vout
** GLOBAL gnd
Rresnwell@0 net@14 gnd 10k
XSingleCe@2 net@11 b3 net@19 Lab_1_DAC__SingleCell
XSingleCe@3 net@8 b2 net@11 Lab_1_DAC__SingleCell
XSingleCe@4 net@13 b1 net@8 Lab_1_DAC__SingleCell
XSingleCe@5 net@14 b0 net@13 Lab_1_DAC__SingleCell
XSingleCe@6 net@19 b4 vout Lab_1_DAC__SingleCell
.ENDS Lab_1_DAC__5BitDAC

.global gnd

*** TOP LEVEL CELL: 5BitDac_sim_digital{sch}
X_5BitDAC@0 net@0 b1 b2 b3 b4 vout Lab_1_DAC__5BitDAC

* Spice Code nodes in cell cell '5BitDac_sim_digital{sch}'
* Digital Input: 10000
Vb4 b4 0 DC 2V
Vb3 b3 0 DC 0V
Vb2 b2 0 DC 0V
Vb1 b1 0 DC 0V
Vb0 b0 0 DC 0V
.op
.END
